module testbench_lab4t1();
 logic a00;
 logic b00;
 logic a11;
 logic b11;
 logic R1;logic G1;logic B1;
 lab4ta dsd(
 .a0(a00),.a1(a11),.b0(b00),.b1(b11),.R(R1),.G(G1), .B(B1)
 );
 initial begin
 a00 = 0; a11 = 0; b00 = 0;b11 = 0;
 #10;
 a00 = 0; a11 = 0; b00 = 0;b11 = 1;
 #10;
 a00 = 0; a11 = 0; b00 = 1;b11 = 0;
 #10;
 a00 = 0; a11 = 0; b00 = 1;b11 = 1;
 #10;
 a00 = 0; a11 = 1; b00 = 0;b11 = 0;
 #10;
 a00 = 0; a11 = 1; b00 = 0;b11 = 1;
 #10;
 a00 = 0; a11 = 1; b00 = 1;b11 = 0;
 #10;
 a00 = 0; a11 = 1; b00 = 1;b11 = 1;
 #10;
 a00 = 1; a11 = 0; b00 = 0;b11 = 0;
 #10;
 a00 = 1; a11 = 0; b00 = 0;b11 = 1;
 #10;
 a00 = 1; a11 = 0; b00 = 1;b11 = 0;
 #10;
 a00 = 1; a11 = 0; b00 = 1;b11 = 1;
 #10;
 a00 = 1; a11 = 1; b00 = 0;b11 = 0;
 #10;
 a00 = 1; a11 = 1; b00 = 0;b11 = 1;
 #10;
 a00 = 1; a11 = 1; b00 = 1;b11 = 0;
 #10;
 a00 = 1; a11 = 1; b00 = 1;b11 = 1;
 #10;
 $stop;
 end 
 endmodule